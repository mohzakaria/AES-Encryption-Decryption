module Cipher_tb;
reg [127:0] in1;
wire [127:0] out1;
reg [127:0] key1;

reg [127:0] in2;
wire [127:0] out2;
reg [191:0] key2;

reg [127:0] in3;
wire [127:0] out3;
reg [255:0] key3;

Cipher a(in1,key1,out1);



initial begin
$monitor("in128= %h, key128= %h ,out128= %h",in1,key1,out1);
in1=128'h00112233445566778899aabbccddeeff;
key1=128'h000102030405060708090a0b0c0d0e0f;
//key=00000000000000010000001000000011000001000000010100000110000001110000100000001001000010100000101100001100000011010000111000001111
//output =69c4e0d86a7b0430d8cdb78070b4c55a
//output binary:01101001110001001110000011011000011010100111101100000100001100001101100011001101101101111000000001110000101101001100010101011010
#10;
end

endmodule
