module SBoxReverse(inputByte,outputByte);
input [7:0] inputByte;
output reg [7:0] outputByte;

always @(*) begin
		case(inputByte)
            8'h63: outputByte= 8'h00;
            8'h7c: outputByte= 8'h01;
            8'h77: outputByte= 8'h02;
            8'h7b: outputByte= 8'h03;
            8'hf2: outputByte= 8'h04;
            8'h6b: outputByte= 8'h05;
            8'h6f: outputByte= 8'h06;
            8'hc5: outputByte= 8'h07;
            8'h30: outputByte=8'h08;
            8'h01: outputByte=8'h09;
            8'h67: outputByte=8'h0a;
            8'h2b: outputByte=8'h0b;
            8'hfe: outputByte=8'h0c;
            8'hd7: outputByte=8'h0d;
            8'hab: outputByte=8'h0e;
            8'h76: outputByte=8'h0f;
            8'hca: outputByte=8'h10;
            8'h82: outputByte=8'h11;
            8'hc9: outputByte=8'h12;
            8'h7d: outputByte=8'h13;
            8'hfa: outputByte=8'h14;
            8'h59: outputByte=8'h15;
            8'h47: outputByte=8'h16; 
            8'hf0: outputByte= 8'h17;
            8'had: outputByte=8'h18;
            8'hd4: outputByte=8'h19;
            8'ha2: outputByte=8'h1a;
            8'haf: outputByte=8'h1b;
            8'h9c: outputByte=8'h1c;
            8'ha4: outputByte=8'h1d;
            8'h72: outputByte=8'h1e;
            8'hc0: outputByte=8'h1f;
            8'hb7: outputByte=8'h20;
            8'hfd: outputByte=8'h21;
            8'h93: outputByte=8'h22;
            8'h26: outputByte=8'h23;
            8'h36: outputByte=8'h24;
            8'h3f: outputByte=8'h25;
            8'hf7: outputByte=8'h26;
            8'hcc: outputByte=8'h27;
            8'h34: outputByte=8'h28;
            8'ha5: outputByte=8'h29;
            8'he5: outputByte=8'h2a;
            8'hf1: outputByte=8'h2b;
            8'h71: outputByte=8'h2c;
            8'hd8: outputByte=8'h2d;
            8'h31: outputByte=8'h2e;
            8'h15: outputByte=8'h2f;
            8'h04: outputByte=8'h30;
            8'hc7: outputByte=8'h31;
            8'h23: outputByte=8'h32;
            8'hc3: outputByte=8'h33;
            8'h18: outputByte=8'h34;
            8'h96: outputByte=8'h35;
            8'h05: outputByte=8'h36;
            8'h9a: outputByte=8'h37;
            8'h07: outputByte=8'h38;
            8'h12: outputByte=8'h39;
            8'h80: outputByte=8'h3a;
            8'he2: outputByte=8'h3b;
            8'heb: outputByte=8'h3c;
            8'h27: outputByte=8'h3d;
            8'hb2: outputByte=8'h3e;
            8'h75: outputByte=8'h3f;
            8'h09: outputByte=8'h40;
            8'h83: outputByte=8'h41;
            8'h2c: outputByte=8'h42;
            8'h1a: outputByte=8'h43;
            8'h1b: outputByte=8'h44;
            8'h6e: outputByte=8'h45;
            8'h5a: outputByte=8'h46;
            8'ha0: outputByte=8'h47;
            8'h52: outputByte=8'h48;
            8'h3b: outputByte=8'h49;
            8'hd6: outputByte=8'h4a;
            8'hb3: outputByte=8'h4b;
            8'h29: outputByte=8'h4c;
            8'he3: outputByte=8'h4d;
            8'h2f: outputByte=8'h4e;
            8'h84: outputByte=8'h4f;
            8'h53: outputByte=8'h50;
            8'hd1: outputByte=8'h51;
            8'h00: outputByte=8'h52;
            8'hed: outputByte=8'h53;
            8'h20: outputByte=8'h54;
            8'hfc: outputByte=8'h55;
            8'hb1: outputByte=8'h56;
            8'h5b: outputByte=8'h57;
            8'h6a: outputByte=8'h58;
            8'hcb: outputByte=8'h59;
            8'hbe: outputByte=8'h5a;
            8'h39: outputByte=8'h5b;
            8'h4a: outputByte=8'h5c;
            8'h4c: outputByte=8'h5d;
            8'h58: outputByte=8'h5e;
            8'hcf: outputByte=8'h5f;
            8'hd0: outputByte=8'h60;
            8'hef: outputByte=8'h61;
            8'haa: outputByte=8'h62;
            8'hfb: outputByte=8'h63;
            8'h43: outputByte=8'h64;
            8'h4d: outputByte=8'h65;
            8'h33: outputByte=8'h66;
            8'h85: outputByte=8'h67;
            8'h45: outputByte=8'h68;
            8'hf9: outputByte=8'h69;
            8'h02: outputByte=8'h6a;
            8'h7f: outputByte=8'h6b;
            8'h50: outputByte=8'h6c;
            8'h3c: outputByte=8'h6d;
            8'h9f: outputByte=8'h6e;
            8'ha8: outputByte=8'h6f;
            8'h51: outputByte=8'h70;
            8'ha3: outputByte=8'h71;
            8'h40: outputByte=8'h72;
            8'h8f: outputByte=8'h73;
            8'h92: outputByte=8'h74;
            8'h9d: outputByte=8'h75;
            8'h38: outputByte=8'h76;
            8'hf5: outputByte=8'h77;
            8'hbc: outputByte=8'h78;
            8'hb6: outputByte=8'h79;
            8'hda: outputByte=8'h7a;
            8'h21: outputByte=8'h7b;
            8'h10: outputByte=8'h7c;
            8'hff: outputByte=8'h7d;
            8'hf3: outputByte=8'h7e;
            8'hd2: outputByte=8'h7f;
            8'hcd: outputByte=8'h80;
            8'h0c: outputByte=8'h81;
            8'h13: outputByte=8'h82;
            8'hec: outputByte=8'h83;
            8'h5f: outputByte=8'h84;
            8'h97: outputByte=8'h85;
            8'h44: outputByte=8'h86;
            8'h17: outputByte=8'h87;
            8'hc4: outputByte=8'h88;
            8'ha7: outputByte=8'h89;
            8'h7e: outputByte=8'h8a;
            8'h3d: outputByte=8'h8b;
            8'h64: outputByte=8'h8c;
            8'h5d: outputByte=8'h8d;
            8'h19: outputByte=8'h8e;
            8'h73: outputByte=8'h8f;
            8'h60: outputByte=8'h90;
            8'h81: outputByte=8'h91;
            8'h4f: outputByte=8'h92;
            8'hdc: outputByte=8'h93;
            8'h22: outputByte=8'h94;
            8'h2a: outputByte=8'h95;
            8'h90: outputByte=8'h96;
            8'h88: outputByte=8'h97;
            8'h46: outputByte=8'h98;
            8'hee: outputByte=8'h99;
            8'hb8: outputByte=8'h9a;
            8'h14: outputByte=8'h9b;
            8'hde: outputByte=8'h9c;
            8'h5e: outputByte=8'h9d;
            8'h0b: outputByte=8'h9e;
            8'hdb: outputByte=8'h9f;
            8'he0: outputByte=8'ha0;
            8'h32: outputByte=8'ha1;
            8'h3a: outputByte=8'ha2;
            8'h0a: outputByte=8'ha3;
            8'h49: outputByte=8'ha4;
            8'h06: outputByte=8'ha5;
            8'h24: outputByte=8'ha6;
            8'h5c: outputByte=8'ha7;
            8'hc2: outputByte=8'ha8;
            8'hd3: outputByte=8'ha9;
            8'hac: outputByte=8'haa;
            8'h62: outputByte=8'hab;
            8'h91: outputByte=8'hac;
            8'h95: outputByte=8'had;
            8'he4: outputByte=8'hae;
            8'h79: outputByte=8'haf;
            8'he7: outputByte=8'hb0;
            8'hc8: outputByte=8'hb1;
            8'h37: outputByte=8'hb2;
            8'h6d: outputByte=8'hb3;
            8'h8d: outputByte=8'hb4;
            8'hd5: outputByte=8'hb5;
            8'h4e: outputByte=8'hb6;
            8'ha9: outputByte=8'hb7;
            8'h6c: outputByte=8'hb8;
            8'h56: outputByte=8'hb9;
            8'hf4: outputByte=8'hba;
            8'hea: outputByte=8'hbb;
            8'h65: outputByte=8'hbc;
            8'h7a: outputByte=8'hbd;
            8'hae: outputByte=8'hbe;
            8'h08: outputByte=8'hbf;
            8'hba: outputByte=8'hc0;
            8'h78: outputByte=8'hc1;
            8'h25: outputByte=8'hc2;
            8'h2e: outputByte=8'hc3;
            8'h1c: outputByte=8'hc4;
            8'ha6: outputByte=8'hc5;
            8'hb4: outputByte=8'hc6;
            8'hc6: outputByte=8'hc7;
            8'he8: outputByte=8'hc8;
            8'hdd: outputByte=8'hc9;
            8'h74: outputByte=8'hca;
            8'h1f: outputByte=8'hcb;
            8'h4b: outputByte=8'hcc;
            8'hbd: outputByte=8'hcd;
            8'h8b: outputByte=8'hce;
            8'h8a: outputByte=8'hcf;
            8'h70: outputByte=8'hd0;
            8'h3e: outputByte=8'hd1;
            8'hb5: outputByte=8'hd2;
            8'h66: outputByte=8'hd3;
            8'h48: outputByte=8'hd4;
            8'h03: outputByte=8'hd5;
            8'hf6: outputByte=8'hd6;
            8'h0e: outputByte=8'hd7;
            8'h61: outputByte=8'hd8;
            8'h35: outputByte=8'hd9;
            8'h57: outputByte=8'hda;
            8'hb9: outputByte=8'hdb;
            8'h86: outputByte=8'hdc;
            8'hc1: outputByte=8'hdd;
            8'h1d: outputByte=8'hde;
            8'h9e: outputByte=8'hdf;
            8'he1: outputByte=8'he0;
            8'hf8: outputByte=8'he1;
            8'h98: outputByte=8'he2;
            8'h11: outputByte=8'he3;
            8'h69: outputByte=8'he4;
            8'hd9: outputByte=8'he5;
            8'h8e: outputByte=8'he6;
            8'h94: outputByte=8'he7;
            8'h9b: outputByte=8'he8;
            8'h1e: outputByte=8'he9;
            8'h87: outputByte=8'hea;
            8'he9: outputByte=8'heb;
            8'hce: outputByte=8'hec;
            8'h55: outputByte=8'hed;
            8'h28: outputByte=8'hee;
            8'hdf: outputByte=8'hef;
            8'h8c: outputByte=8'hf0;
            8'ha1: outputByte=8'hf1;
            8'h89: outputByte=8'hf2;
            8'h0d: outputByte=8'hf3;
            8'hbf: outputByte=8'hf4;
            8'he6: outputByte=8'hf5;
            8'h42: outputByte=8'hf6;
            8'h68: outputByte=8'hf7;
            8'h41: outputByte=8'hf8;
            8'h99: outputByte=8'hf9;
            8'h2d: outputByte=8'hfa;
            8'h0f: outputByte=8'hfb;
            8'hb0: outputByte=8'hfc;
            8'h54: outputByte=8'hfd;
            8'hbb: outputByte=8'hfe;
            8'h16: outputByte=8'hff;
			default: 
			outputByte = 8'h00;
		endcase
	end
endmodule 