module ProjectLogic2(inputState,outputState);
input [127:0] inputState;
output [127:0] outputState;



endmodule 

